library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use work.ML_types.all;
use work.CNN_W_cnn1.all;
use work.CNN_W_cnn2.all;
use work.CNN_W_fc.all;

entity tb_CNN is
end entity;

-- an example of a test bench
architecture test of tb_CNN is

    component CNN is
        port (
            CLK  : in std_logic;
            RSTn : in std_logic;
            I : in tensor2D (0 to 28) (0 to 28) (7 downto 0);
            O : out std_logic_vector(9 downto 0);
            DONE : out std_logic
        );
    end component;

    signal CLK  : std_logic := '0';
    signal RSTn : std_logic := '0';
    
    -- number 7
    signal I : tensor2D (0 to 28) (0 to 28) (7 downto 0) := (
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"d4", x"39", x"1f", x"17", x"bc", x"a4", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"5e", x"7e", x"7e", x"7e", x"7e", x"71", x"46", x"46", x"46", x"46", x"46", x"46", x"46", x"46", x"2a", x"b4", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"c3", x"f2", x"c8", x"f2", x"23", x"63", x"7e", x"61", x"7e", x"7e", x"7e", x"7a", x"65", x"7e", x"7e", x"0c", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"91", x"c2", x"8e", x"c3", x"c3", x"c3", x"bb", x"95", x"6c", x"7e", x"ea", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"d3", x"7d", x"51", x"92", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"96", x"69", x"7f", x"d3", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"01", x"7e", x"6e", x"ac", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"bb", x"79", x"7e", x"be", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"05", x"7e", x"3b", x"85", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"89", x"4d", x"78", x"ba", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"fe", x"7e", x"36", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"cb", x"7b", x"70", x"b9", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"93", x"5d", x"7e", x"26", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"83", x"4b", x"7e", x"5b", x"a3", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"a6", x"7e", x"7e", x"cd", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"9f", x"60", x"7e", x"f3", x"81", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"05", x"7e", x"7e", x"b4", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"bd", x"72", x"7e", x"7e", x"b4", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"f9", x"7e", x"7e", x"5b", x"a8", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"f9", x"7e", x"4f", x"92", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
        (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80")
    );

    -- -- number 2
    -- signal I : tensor2D (0 to 28) (0 to 28) (7 downto 0) := (
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"f4", x"fd", x"2b", x"7f", x"7f", x"16", x"dd", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"29", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"5a", x"9e", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"29", x"7d", x"7d", x"7d", x"55", x"0e", x"30", x"7d", x"7d", x"fa", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"b4", x"7a", x"7d", x"52", x"a0", x"8c", x"80", x"86", x"4e", x"7d", x"0c", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"cd", x"7b", x"52", x"99", x"80", x"80", x"80", x"fa", x"78", x"7d", x"c1", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"9f", x"92", x"80", x"80", x"80", x"80", x"51", x"7d", x"7d", x"c1", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"f5", x"77", x"7d", x"46", x"8a", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"cc", x"77", x"7d", x"67", x"bf", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"7d", x"7d", x"10", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"30", x"76", x"7d", x"1f", x"8c", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"99", x"6a", x"7d", x"69", x"a3", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"46", x"7d", x"7d", x"0d", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"ce", x"78", x"7d", x"3d", x"8c", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"93", x"48", x"7d", x"7d", x"0d", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"06", x"7d", x"7d", x"2d", x"8c", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"78", x"7d", x"7d", x"99", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"78", x"7d", x"7d", x"ab", x"94", x"94", x"94", x"94", x"85", x"80", x"85", x"94", x"94", x"a5", x"16", x"16", x"16", x"13", x"8a", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"78", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"28", x"0f", x"26", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"fb", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"2e", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"79", x"77", x"77", x"29", x"f5", x"f5", x"b9", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"f6", x"fb", x"fb", x"fb", x"26", x"7d", x"7d", x"7d", x"1b", x"fb", x"fb", x"a9", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"),
    --     (x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80")
    -- );

    signal O : std_logic_vector(9 downto 0);
    signal DONE : std_logic;

    begin

        CNN_dut: CNN port map (CLK => CLK, RSTn => RSTn, I => I, O => O, DONE => DONE);

        -- clock process
        process
        begin
            while true loop
                clk <= '0';
                wait for 5 ns;
                clk <= '1';
                wait for 5 ns;
            end loop;
        end process;

        -- reset
        RSTn <= '0', '1' after 20 ns;

end architecture;
